* NGSPICE file created from sky130_ef_ip__template.ext - technology: sky130A

.subckt sky130_ef_ip__template A Y VPWR VGND
X0 Y.t0 A.t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 Y.t1 A.t1 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 A.n0 A.t1 396.195
R1 A.n0 A.t0 381.74
R2 A A.n0 0.8755
R3 VGND.n7 VGND.n3 2126.44
R4 VGND.n4 VGND.n1 2126.44
R5 VGND.n5 VGND.n4 776.759
R6 VGND.n7 VGND.n6 776.759
R7 VGND.n3 VGND.n2 292.5
R8 VGND.n9 VGND.n1 292.5
R9 VGND.n5 VGND.n3 163.206
R10 VGND.n6 VGND.n1 163.206
R11 VGND.n4 VGND.n0 146.25
R12 VGND.n8 VGND.n7 146.25
R13 VGND.n2 VGND.n0 138.166
R14 VGND.n9 VGND.n0 138.166
R15 VGND.n8 VGND.n2 138.166
R16 VGND.n9 VGND.n8 138.166
R17 VGND.n6 VGND.t0 106.847
R18 VGND.t0 VGND.n5 106.847
R19 VGND.n10 VGND.t1 84.1063
R20 VGND.n10 VGND.n9 1.93237
R21 VGND VGND.n10 0.227062
R22 Y.n0 Y.t1 229.275
R23 Y.n0 Y.t0 84.8468
R24 Y Y.n0 0.516125
R25 VPWR.n7 VPWR.n1 1312.94
R26 VPWR.n5 VPWR.n4 1312.94
R27 VPWR.n4 VPWR.n3 237.584
R28 VPWR.n7 VPWR.n6 237.584
R29 VPWR.n10 VPWR.t1 228.589
R30 VPWR.n9 VPWR.n8 140.048
R31 VPWR.n8 VPWR.n2 140.048
R32 VPWR.n2 VPWR.n0 140.048
R33 VPWR.n9 VPWR.n0 140.048
R34 VPWR.n5 VPWR.n2 92.5005
R35 VPWR.n9 VPWR.n1 92.5005
R36 VPWR.n3 VPWR.n1 70.7763
R37 VPWR.n6 VPWR.n5 70.7763
R38 VPWR.n8 VPWR.n7 46.2505
R39 VPWR.n4 VPWR.n0 46.2505
R40 VPWR.n6 VPWR.t0 16.7394
R41 VPWR.n3 VPWR.t0 16.7394
R42 VPWR.n10 VPWR.n9 1.93237
R43 VPWR VPWR.n10 0.227062
C0 Y VPWR 0.34468f
C1 A VPWR 0.246347f
C2 A Y 0.233998f
C3 Y VGND 0.546265f
C4 A VGND 0.432827f
C5 VPWR VGND 1.27866f
.ends

