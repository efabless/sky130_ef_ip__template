* NGSPICE file created from sky130_ef_ip__template.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_D5KUY4 a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_ZUW952 a_n73_n64# a_n33_n161# a_15_n64# w_n211_n284#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n211_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_ef_ip__template A Y VPWR VGND
XXM1 Y VGND A VGND sky130_fd_pr__nfet_01v8_D5KUY4
XXM2 VPWR A Y VPWR sky130_fd_pr__pfet_01v8_ZUW952
.ends

